`define BusOwner 1:0
`define BUS_MASTER_NUM 4
`define BUS_MASTER_0 2'h0
`define BUS_MASTER_1 2'h1
`define BUS_MASTER_2 2'h2
`define BUS_MASTER_3 2'h3

`define BusSlaveIndex 2:0
`define BusSlaveIndexLoc 29:27
`define BUS_SLAVE_INDEX_NUM 3
`define BUS_SLAVE_NUM 8
`define BUS_SLAVE_0 0
`define BUS_SLAVE_1 1
`define BUS_SLAVE_2 2
`define BUS_SLAVE_3 3
`define BUS_SLAVE_4 4
`define BUS_SLAVE_5 5
`define BUS_SLAVE_6 6
`define BUS_SLAVE_7 7
