`define ROM_SIZE 8192
`define ROM_DEPTH 2048
`define ROM_ADDR_W 11
`define RomAddr 10:0
`define RomAddrLoc 10:0