`ifndef __GLOBAL_CONFIG_VH__
`define __GLOBAL_CONFIG_VH__

`define RST_EDGE negedge
`define RST_ENABLE 1'b0
`define RST_DISABLE 1'b1

`define MEM_ENABLE 1'b1
`define MEM_DISABLE 1'b0

`endif