`define ISA_NOP 32'h0
`define ISA_OP_W 6
`define IsaOpBus 5:0