// 16384 = 4096 * 4 (there is 4 bytes in a word since the cpu is 32-bit)
`define SPM_SIZE 16384
`define SPM_DEPTH 4096
`define SPM_ADDR_W 12

`define SpmAddrBus 11:0
`define SpmAddrLoc 11:0
